// JTAG TAP Controller Testbench
// Designer: Copilot
//
// Unit test for IEEE 1149.1 compliant TAP controller

`timescale 1ns/1ps

module test_tap_controller;

    // Test parameters
    localparam real TCK_PERIOD_NS = 100.0;  // 10 MHz TCK (100ns period)
    localparam int  TEST_TIMEOUT_CYCLES = 10000;

    // JTAG Signals
    logic TCK;
    logic TMS;
    logic TDI;
    logic TDO;
    logic TRST_n;

    // IJTAG Interface
    logic ijtag_select;
    logic ijtag_capture;
    logic ijtag_shift;
    logic ijtag_update;
    logic ijtag_tdi;
    logic ijtag_tdo;

    // Instantiate DUT
    tap_controller dut (
        .TCK           (TCK),
        .TMS           (TMS),
        .TDI           (TDI),
        .TDO           (TDO),
        .TRST_n        (TRST_n),
        .ijtag_select  (ijtag_select),
        .ijtag_capture (ijtag_capture),
        .ijtag_shift   (ijtag_shift),
        .ijtag_update  (ijtag_update),
        .ijtag_tdi     (ijtag_tdi),
        .ijtag_tdo     (ijtag_tdo)
    );

    // TCK generation (10 MHz = 100 ns period)
    initial begin
        TCK = 0;
        forever #(TCK_PERIOD_NS/2) TCK = ~TCK;
    end

    // Test stimulus
    initial begin
        // Initialize signals
        TMS     = 1;
        TDI     = 0;
        TRST_n  = 0;
        ijtag_tdo = 0;

        // Generate waveform dump
        $dumpfile("test_tap_controller.vcd");
        $dumpvars(0, test_tap_controller);

        $display("=== JTAG TAP Controller Test Started ===");
        $display("TCK Period: %.1f ns (%.1f MHz)", TCK_PERIOD_NS, 1000.0/TCK_PERIOD_NS);

        // Release reset
        #(TCK_PERIOD_NS * 2);
        TRST_n = 1;
        #(TCK_PERIOD_NS * 2);

        // Test 1: TAP Reset and IDLE
        $display("\n[Test 1] Testing TAP Reset and Run-Test-Idle");
        tap_reset();
        check_state_reset();
        goto_idle();
        $display("[Test 1] PASS - TAP in Run-Test-Idle state");

        // Test 2: Instruction Register Scan
        $display("\n[Test 2] Testing Instruction Register Scan");
        tap_reset();
        goto_idle();
        
        // Load IDCODE instruction
        shift_ir(4'h1);
        $display("[Test 2] Loaded IDCODE instruction");
        
        // Load BYPASS instruction
        shift_ir(4'h0);
        $display("[Test 2] Loaded BYPASS instruction");
        
        // Load TCP_CTRL instruction
        shift_ir(4'h8);
        $display("[Test 2] Loaded TCP_CTRL instruction");
        
        $display("[Test 2] PASS - Instruction register operations");

        // Test 3: BYPASS Data Register
        $display("\n[Test 3] Testing BYPASS Data Register");
        tap_reset();
        goto_idle();
        shift_ir(4'h0);  // BYPASS instruction
        
        // Shift through BYPASS (1 bit)
        goto_shift_dr();
        @(posedge TCK);
        TDI = 1;
        TMS = 0;  // Stay in SHIFT-DR
        @(negedge TCK);
        // TDO should still be 0 (previous BYPASS value)
        if (TDO == 0) begin
            $display("[Test 3] First shift: TDO=0 (previous value) - correct");
        end else begin
            $display("[Test 3] FAIL - Expected TDO=0, got TDO=%b", TDO);
        end
        @(posedge TCK);
        TDI = 0;
        TMS = 1;  // Exit SHIFT-DR
        @(negedge TCK);
        // Now TDO should be 1 (the value we shifted in)
        if (TDO == 1) begin
            $display("[Test 3] PASS - BYPASS shifted correctly, TDO=1");
        end else begin
            $display("[Test 3] FAIL - BYPASS expected TDO=1, got TDO=%b", TDO);
        end
        goto_idle();

        // Test 4: IDCODE Data Register
        $display("\n[Test 4] Testing IDCODE Data Register");
        tap_reset();
        // After reset, IDCODE should be selected by default
        goto_shift_dr();
        
        // Shift out 32 bits of IDCODE
        logic [31:0] idcode_read;
        for (int i = 0; i < 32; i++) begin
            @(posedge TCK);
            TDI = 0;
            TMS = (i == 31) ? 1 : 0;  // Exit on last bit
            @(negedge TCK);
            idcode_read[i] = TDO;
        end
        
        // Expected IDCODE: {4'h1, 16'hCAFE, 11'h05F, 1'b1}
        logic [31:0] expected_idcode = {4'h1, 16'hCAFE, 11'h05F, 1'b1};
        if (idcode_read == expected_idcode) begin
            $display("[Test 4] PASS - IDCODE read: 0x%08h", idcode_read);
        end else begin
            $display("[Test 4] FAIL - Expected 0x%08h, got 0x%08h", expected_idcode, idcode_read);
        end
        goto_idle();

        // Test 5: TCP_CTRL Write and Read
        $display("\n[Test 5] Testing TCP_CTRL Register");
        tap_reset();
        goto_idle();
        shift_ir(4'h8);  // TCP_CTRL instruction
        
        // Write test pattern to TCP_CTRL
        logic [31:0] test_pattern = 32'hA5A5_5A5A;
        shift_dr_32(test_pattern);
        
        // Read back TCP_CTRL
        logic [31:0] readback;
        shift_dr_32_read(readback);
        
        if (readback == test_pattern) begin
            $display("[Test 5] PASS - TCP_CTRL write/read: 0x%08h", readback);
        end else begin
            $display("[Test 5] FAIL - Expected 0x%08h, got 0x%08h", test_pattern, readback);
        end

        // Test 6: TCP_STATUS Read (Read-only register)
        $display("\n[Test 6] Testing TCP_STATUS Register");
        tap_reset();
        goto_idle();
        shift_ir(4'h9);  // TCP_STATUS instruction
        
        // Read TCP_STATUS
        logic [31:0] status;
        shift_dr_32_read(status);
        $display("[Test 6] TCP_STATUS read: 0x%08h (expected 0xDEADBEEF)", status);
        
        if (status == 32'hDEAD_BEEF) begin
            $display("[Test 6] PASS - TCP_STATUS read correctly");
        end else begin
            $display("[Test 6] FAIL - Expected 0xDEADBEEF, got 0x%08h", status);
        end

        // Test 7: IJTAG_ACCESS Instruction
        $display("\n[Test 7] Testing IJTAG_ACCESS Instruction");
        tap_reset();
        goto_idle();
        shift_ir(4'hA);  // IJTAG_ACCESS instruction
        
        // Check IJTAG interface signals
        goto_capture_dr();
        @(posedge TCK);
        if (ijtag_select && ijtag_capture) begin
            $display("[Test 7] IJTAG select and capture asserted");
        end else begin
            $display("[Test 7] FAIL - IJTAG signals not asserted (select=%b, capture=%b)", 
                     ijtag_select, ijtag_capture);
        end
        
        goto_shift_dr();
        @(posedge TCK);
        if (ijtag_select && ijtag_shift) begin
            $display("[Test 7] PASS - IJTAG shift asserted");
        end else begin
            $display("[Test 7] FAIL - IJTAG shift not asserted");
        end
        goto_idle();

        // Test 8: State Transitions
        $display("\n[Test 8] Testing Complete State Machine Transitions");
        tap_reset();
        test_all_states();
        $display("[Test 8] PASS - All state transitions verified");

        // Test 9: TCK Frequency Verification (max 10 MHz)
        $display("\n[Test 9] Verifying TCK Frequency");
        if (TCK_PERIOD_NS >= 100.0) begin
            $display("[Test 9] PASS - TCK period %.1f ns (%.1f MHz) <= 10 MHz", 
                     TCK_PERIOD_NS, 1000.0/TCK_PERIOD_NS);
        end else begin
            $display("[Test 9] FAIL - TCK frequency exceeds 10 MHz");
        end

        // Test 10: Multiple Instruction Switches
        $display("\n[Test 10] Testing Multiple Instruction Switches");
        tap_reset();
        goto_idle();
        
        shift_ir(4'h1);  // IDCODE
        shift_ir(4'h0);  // BYPASS
        shift_ir(4'h8);  // TCP_CTRL
        shift_ir(4'h9);  // TCP_STATUS
        shift_ir(4'hA);  // IJTAG_ACCESS
        
        $display("[Test 10] PASS - Multiple instruction switches completed");

        $display("\n=== All Tests Completed Successfully ===");
        #(TCK_PERIOD_NS * 10);
        $finish;
    end

    // Helper Tasks

    // Reset TAP to TEST-LOGIC-RESET state
    task tap_reset();
        @(posedge TCK);
        TMS = 1;
        repeat(5) @(posedge TCK);  // 5 TMS=1 transitions guarantee reset
        $display("  TAP reset to TEST-LOGIC-RESET");
    endtask

    // Check if in TEST-LOGIC-RESET state
    task check_state_reset();
        if (dut.tap_state == dut.TEST_LOGIC_RESET) begin
            $display("  Confirmed in TEST-LOGIC-RESET state");
        end else begin
            $display("  ERROR: Not in TEST-LOGIC-RESET state");
        end
    endtask

    // Go to RUN-TEST-IDLE state
    task goto_idle();
        @(posedge TCK);
        TMS = 0;  // From TEST-LOGIC-RESET to RUN-TEST-IDLE (or stay in RUN-TEST-IDLE)
        @(posedge TCK);
    endtask

    // Go to SHIFT-IR state
    task goto_shift_ir();
        @(posedge TCK);
        TMS = 1;  // SELECT-DR-SCAN
        @(posedge TCK);
        TMS = 1;  // SELECT-IR-SCAN
        @(posedge TCK);
        TMS = 0;  // CAPTURE-IR
        @(posedge TCK);
        TMS = 0;  // SHIFT-IR
        @(posedge TCK);
    endtask

    // Go to SHIFT-DR state
    task goto_shift_dr();
        @(posedge TCK);
        TMS = 1;  // SELECT-DR-SCAN
        @(posedge TCK);
        TMS = 0;  // CAPTURE-DR
        @(posedge TCK);
        TMS = 0;  // SHIFT-DR
        @(posedge TCK);
    endtask

    // Go to CAPTURE-DR state
    task goto_capture_dr();
        @(posedge TCK);
        TMS = 1;  // SELECT-DR-SCAN
        @(posedge TCK);
        TMS = 0;  // CAPTURE-DR
        @(posedge TCK);
    endtask

    // Shift Instruction Register (4 bits)
    task shift_ir(input logic [3:0] instruction);
        goto_shift_ir();
        
        for (int i = 0; i < 4; i++) begin
            @(posedge TCK);
            TDI = instruction[i];
            TMS = (i == 3) ? 1 : 0;  // Exit on last bit
        end
        
        // Update-IR
        @(posedge TCK);
        TMS = 1;  // Go to UPDATE-IR
        @(posedge TCK);
        TMS = 0;  // Go to RUN-TEST-IDLE
        @(posedge TCK);
    endtask

    // Shift Data Register (32 bits) - Write
    task shift_dr_32(input logic [31:0] data);
        goto_shift_dr();
        
        for (int i = 0; i < 32; i++) begin
            @(posedge TCK);
            TDI = data[i];
            TMS = (i == 31) ? 1 : 0;  // Exit on last bit
        end
        
        // Update-DR
        @(posedge TCK);
        TMS = 1;  // Go to UPDATE-DR
        @(posedge TCK);
        TMS = 0;  // Go to RUN-TEST-IDLE
        @(posedge TCK);
    endtask

    // Shift Data Register (32 bits) - Read
    task shift_dr_32_read(output logic [31:0] result);
        goto_shift_dr();
        
        for (int i = 0; i < 32; i++) begin
            @(posedge TCK);
            TDI = 0;
            TMS = (i == 31) ? 1 : 0;  // Exit on last bit
            @(negedge TCK);
            result[i] = TDO;
        end
        
        // Update-DR
        @(posedge TCK);
        TMS = 1;  // Go to UPDATE-DR
        @(posedge TCK);
        TMS = 0;  // Go to RUN-TEST-IDLE
        @(posedge TCK);
    endtask

    // Test all state transitions
    task test_all_states();
        // Test DR path
        TMS = 1; @(posedge TCK);  // SELECT-DR-SCAN
        TMS = 0; @(posedge TCK);  // CAPTURE-DR
        TMS = 0; @(posedge TCK);  // SHIFT-DR
        TMS = 1; @(posedge TCK);  // EXIT1-DR
        TMS = 0; @(posedge TCK);  // PAUSE-DR
        TMS = 1; @(posedge TCK);  // EXIT2-DR
        TMS = 0; @(posedge TCK);  // SHIFT-DR
        TMS = 1; @(posedge TCK);  // EXIT1-DR
        TMS = 1; @(posedge TCK);  // UPDATE-DR
        TMS = 0; @(posedge TCK);  // RUN-TEST-IDLE
        
        // Test IR path
        TMS = 1; @(posedge TCK);  // SELECT-DR-SCAN
        TMS = 1; @(posedge TCK);  // SELECT-IR-SCAN
        TMS = 0; @(posedge TCK);  // CAPTURE-IR
        TMS = 0; @(posedge TCK);  // SHIFT-IR
        TMS = 1; @(posedge TCK);  // EXIT1-IR
        TMS = 0; @(posedge TCK);  // PAUSE-IR
        TMS = 1; @(posedge TCK);  // EXIT2-IR
        TMS = 0; @(posedge TCK);  // SHIFT-IR
        TMS = 1; @(posedge TCK);  // EXIT1-IR
        TMS = 1; @(posedge TCK);  // UPDATE-IR
        TMS = 0; @(posedge TCK);  // RUN-TEST-IDLE
        
        $display("  Completed full state machine traversal");
    endtask

    // Timeout watchdog
    initial begin
        #(TCK_PERIOD_NS * TEST_TIMEOUT_CYCLES);
        $display("ERROR: Test timeout!");
        $error("Simulation exceeded maximum time limit");
        $finish;
    end

endmodule
